module data_path #(

)(

);

endmodule