module RISCV32I(
    output logic [31:0]
);


    logic branch_ex


endmodule